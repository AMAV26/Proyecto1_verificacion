//Agente-Generador

class agente (#parameter pkgsize = 16, parameter drvrs=4;)
    